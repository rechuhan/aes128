
`include "aes128_base_test.sv"
`include "aes128_simple_test/aes128_simple_test.sv"



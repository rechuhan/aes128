
`include "aes128_base_test.sv"
//`include "aes128_simple_test/aes128_simple_test.sv"
`include "aes128_direct_test/aes128_direct_test.sv"
`include "aes128_rand_test/aes128_rand_test.sv"


`ifndef __TB_PKG_SV__
`define __TB_PKG_SV__

package tb_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import crypto_dpi_pkg::*;
import aes128_pkg::*;
`include "virtual_sequencer.sv"
`include "tb.sv"

endpackage

`endif

